`ifndef APB_PACKAGE_SVH
`define APB_PACKAGE_SVH

package apb_package;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    
    `include "apb_config.sv"
    `include "apb_define.svh"
    `include "apb_if.sv"
    `include "apb_seq_item.sv"
    `include "apb_driver_base.sv"
    `include "apb_monitor_base.sv"
    `include "apb_master_driver.sv"
    `include "apb_master_monitor.sv"
    `include "apb_agent_base.sv"
    `include "apb_master_agent.sv"
    `include "apb_slave_agent.sv"
    `include "apb_env_base.sv"
    `include "apb_master_env.sv"
    `include "apb_slave_env.sv"
    
    `include "apb_master_basic_seq.sv"
    `include "apb_master_basic_rw_test.sv"

endpackage

`endif