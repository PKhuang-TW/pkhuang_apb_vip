`ifndef APB_DEFINE_SVH
`define APB_DEFINE_SVH

`define     D_ADDR_WIDTH        32
`define     D_DATA_WIDTH        16
`define     D_SLV_COUNT         1

`endif