`ifndef APB_PACKAGE_SVH
`define APB_PACKAGE_SVH

package apb_package;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    
    `include "apb_define.svh"
    `include "apb_interface.sv"
    `include "apb_seq_item.sv"
    `include "apb_driver_base.sv"
    `include "apb_monitor_base.sv"
    `include "apb_master_driver.sv"
    `include "apb_master_monitor.sv"
    `include "apb_slave_driver.sv"
    `include "apb_slave_monitor.sv"
    `include "apb_agent_base.sv"
    `include "apb_master_agent.sv"
    `include "apb_slave_agent.sv"
    `include "apb_scoreboard.sv"
    `include "apb_coverage.sv"
    `include "apb_env.sv"

    `include "apb_master_seq.sv"
    `include "apb_slave_seq.sv"
    `include "apb_basic_rw_test.sv"

endpackage

`endif