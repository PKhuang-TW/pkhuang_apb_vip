`ifndef APB_DEFINE_SVH
`define APB_DEFINE_SVH

`define     D_ADDR_WIDTH        64
`define     D_DATA_WIDTH        32
`define     D_SLV_COUNT         1

`define     D_MEM_SIZE          256

typedef enum { MST, SLV }       apb_role_e;

`endif